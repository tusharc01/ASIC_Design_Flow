/home/nitrkl9/Documents/lock_files/PhysicalDesign/Dependency_Files_GUI/LEF_Files/tsl18fs120_scl.lef